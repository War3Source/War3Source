-- File:
-- Author:
-- Date:
-- Revision:
-- Description:

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.numeric_bit.all;
use std.textio.all;
use ieee.std_logic_textio.all;


-- ENTITY DECLARATION ------------------------------------------------------------------------------
entity _H_ is
      -- generic / port / local declatations
end entity _H_;


-- ARCHITECTURE DECLARATION ------------------------------------------------------------------------
architecture _H_ of _H_ is
     -- local declarations (use function type file component constant signal procedure subtype alias)
begin
     
end architecture _H_;

